Begin3
Language:    SV, 850, Swedish
Description: N�tverksbaserad pakethanterare
Keywords:    fdnpkg16,fdnpkg,uppdatering,paket
End
