Begin3
Language:    SV, 850, Swedish
Description: N�tverksbaserad pakethanterare
Keywords:    fdnpkg,uppdatering,paket
End
